module gNot (input a, output not_a) begin

	assign not_a = !a;

end