module new_gNot (input a, output not_a);

	assign not_a = !a;

endmodule